`timescale 1ns/1ps

// module seg7 (CA, CB, CC, CD, CE, CF, CG, DP, AN);